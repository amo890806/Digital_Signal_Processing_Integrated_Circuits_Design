`define ORDER 23
`define DATA_WIDTH 16
`define ROM_INPUT_MEM_SIZE 40000
`define ROM_OUTPUT_MEM_SIZE 40023
`define FIFO_SIZE 25